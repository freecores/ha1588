`timescale 1ns/1ns

module reg (
);

endmodule
