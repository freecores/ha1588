`timescale 1ns/1ns

module top (
);

endmodule
